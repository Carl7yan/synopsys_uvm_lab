package packet_seq_lib_pkg;
  import uvm_pkg::*;

  class packet extends uvm_sequence_item;
    rand bit[3:0] sa, da;
    rand bit[7:0] payload[$];

    `uvm_object_utils_begin(packet)
      `uvm_field_int(sa, UVM_ALL_ON | UVM_NOCOMPARE)
      `uvm_field_int(da, UVM_ALL_ON)
      `uvm_field_queue_int(payload, UVM_ALL_ON)
    `uvm_object_utils_end

    constraint valid {
      payload.size inside {[1:10]};
    }

    function new(string name="packet");
      super.new(name);
      `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH)
    endfunction
  endclass

  class packet_seq_lib extends uvm_sequence_library #(packet);
  `uvm_object_utils(packet_seq_lib)
  `uvm_sequence_library_utils(packet_seq_lib)

    function new(string name = "packet_seq_lib");
      super.new(name);
      `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
      init_sequence_library();
    endfunction
  endclass


endpackage
